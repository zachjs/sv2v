// pattern: unexpected token 'highz1'
module top;
    wire (highz0, highz1) x;
endmodule
