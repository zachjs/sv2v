module top;
    logic y;
    y = 1;
endmodule
