// pattern: Reached EOF while looking for: "\*/"
/*
