// pattern: compiler directives are forbidden inside strings
`"asdf `line`"
