`START
`ifdef DEFINED
`ifndef NOT_DEFINED
    initial $display("Hi");
`endif
`endif
`END
