module top;
    wire x;
    wire [2:0] y;
    assign y = 1'sb1;
endmodule
