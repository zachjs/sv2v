module top;
    wire [1:0] o1;
    Test1 bar(o1);
    wire o2;
    Test2 test2(o2);
    wire o3;
    Test3 test3(o3);
endmodule
