module top;
    real r = 3.14;
    initial $display(r);
endmodule
