module one;
    logic x;
endmodule
