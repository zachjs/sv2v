module top;
`define PRINT(str) initial $display(`"str`");
`PRINT(a)
`PRINT(\\)
endmodule
