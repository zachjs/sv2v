// pattern: unexpected end of input
`define MACRO(a)
`MACRO
