// pattern: could not find class "C"
module top;
    initial $display(C#()::X);
endmodule
