// pattern: unexpected end of input, looking for '>'
`include <foo
