`ifdef FOO
