// pattern: element "yes" has mismatched end label "no"
module top;
    function yes;
        yes = 0;
    endfunction : no
endmodule
