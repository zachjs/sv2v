// pattern: `endif directive outside of an `if/`endif block
`endif
