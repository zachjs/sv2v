// pattern: decl_bare\.sv:3:5: Parse error: declaration missing type information
module top;
    a;
endmodule
