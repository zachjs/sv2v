module top;
    localparam FOO = 1;
    initial $display(FOO);
endmodule
