// pattern: localparam "X" has no default value
module top;
    localparam X;
endmodule
