// pattern: missing expected `endpackage`
package foo;
