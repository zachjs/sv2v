module surprise;
    initial $display("This isn't what you're looking for!");
endmodule
