module top;
    apple a();
    orange o();
endmodule
