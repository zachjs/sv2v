// pattern: const_const\.sv:3:11: Parse error: duplicate const modifier
module top;
    const const logic x = 1'b1;
endmodule
