// pattern: missing expected `endtask`
module top;
    task automatic foo;
        input inp;
endmodule
