`line 1 "asd" 1B
