module Example;
    reg [15:0] t;
    initial begin
        $display(" 0 xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx xxxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 1 0000001xxxxxxxxxxxxxxxxxxxxxxxxxxxxxx 0000001 xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 2 0000111xxxxxxxxxxxxxxxxxxxxxxxxxxxxxx 0000111 xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 3 0011111xxxxxxxxxxxxxxxxxxxxxxxxxxxxxx 0011111 xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 4 1011111xxxxxxxxxxxxxxxxxxxxxxxxxxxxxx 1011111 xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 5 1010111xxxxxxxxxxxxxxxxxxxxxxxxxxxxxx 1010111 xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 6 10101111xxxxxxxxxxxxxxxxxxxxxxxxxxxxx 1010111 1xx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 7 101011101xxxxxxxxxxxxxxxxxxxxxxxxxxxx 1010111 01x xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 8 1010111010xxxxxxxxxxxxxxxxxxxxxxxxxxx 1010111 010 xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display(" 9 1010111001xxxxxxxxxxxxxxxxxxxxxxxxxxx 1010111 001 xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("11 1010111001xx1xxxxxxxxxxxxxxxxxxxxxxxx 1010111 001 xx1 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("12 1010111001x01xxxxxxxxxxxxxxxxxxxxxxxx 1010111 001 x01 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("13 1010111001001xxxxxxxxxxxxxxxxxxxxxxxx 1010111 001 001 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("14 1010111001011xxxxxxxxxxxxxxxxxxxxxxxx 1010111 001 011 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("15 1010111001001xxxxxxxxxxxxxxxxxxxxxxxx 1010111 001 001 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("16 1010111001001x1xxxxxxxxxxxxxxxxxxxxxx 1010111 001 001 x1xxxx x1x xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("17 1010111001001x01xxxxxxxxxxxxxxxxxxxxx 1010111 001 001 x01xxx x01 xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("18 1010111001001001xxxxxxxxxxxxxxxxxxxxx 1010111 001 001 001xxx 001 xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("19 1010111001001010xxxxxxxxxxxxxxxxxxxxx 1010111 001 001 010xxx 010 xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("20 1010111001001001xxxxxxxxxxxxxxxxxxxxx 1010111 001 001 001xxx 001 xxx xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("21 1010111001001111111xxxxxxxxxxxxxxxxxx 1010111 001 001 111111 111 111 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("22 1010111001001111011xxxxxxxxxxxxxxxxxx 1010111 001 001 111011 111 011 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("23 1010111001001111000xxxxxxxxxxxxxxxxxx 1010111 001 001 111000 111 000 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("24 1010111001001010011xxxxxxxxxxxxxxxxxx 1010111 001 001 010011 010 011 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("25 1010111001001101011xxxxxxxxxxxxxxxxxx 1010111 001 001 101011 101 011 xxxxxx xxx xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("26 1010111001001101011xxxx1xxxxxxxxxxxxx 1010111 001 001 101011 101 011 xxxx1x x1x xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("27 1010111001001101011xxxx01xxxxxxxxxxxx 1010111 001 001 101011 101 011 xxxx01 x01 xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("28 1010111001001101011xxx001xxxxxxxxxxxx 1010111 001 001 101011 101 011 xxx001 001 xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("29 1010111001001101011xxx010xxxxxxxxxxxx 1010111 001 001 101011 101 011 xxx010 010 xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("30 1010111001001101011xxx001xxxxxxxxxxxx 1010111 001 001 101011 101 011 xxx001 001 xxx xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("31 1010111001001101011111111xxxxxxxxxxxx 1010111 001 001 101011 101 011 111111 111 111 xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("32 1010111001001101011011111xxxxxxxxxxxx 1010111 001 001 101011 101 011 011111 111 011 xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("33 1010111001001101011000111xxxxxxxxxxxx 1010111 001 001 101011 101 011 000111 111 000 xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("34 1010111001001101011010011xxxxxxxxxxxx 1010111 001 001 101011 101 011 010011 011 010 xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("35 1010111001001101011101011xxxxxxxxxxxx 1010111 001 001 101011 101 011 101011 011 101 xxxxxx xxx xxx xxxxxx xxx xxx");
        $display("36 1010111001001101011101011x1xxxxxxxxxx 1010111 001 001 101011 101 011 101011 011 101 x1xxxx x1x xxx xxxxxx xxx xxx");
        $display("37 101011100100110101110101101xxxxxxxxxx 1010111 001 001 101011 101 011 101011 011 101 01xxxx 01x xxx xxxxxx xxx xxx");
        $display("38 1010111001001101011101011000xxxxxxxxx 1010111 001 001 101011 101 011 101011 011 101 000xxx 000 xxx xxxxxx xxx xxx");
        $display("39 1010111001001101011101011100xxxxxxxxx 1010111 001 001 101011 101 011 101011 011 101 100xxx 100 xxx xxxxxx xxx xxx");
        $display("40 1010111001001101011101011010xxxxxxxxx 1010111 001 001 101011 101 011 101011 011 101 010xxx 010 xxx xxxxxx xxx xxx");
        $display("41 1010111001001101011101011111111xxxxxx 1010111 001 001 101011 101 011 101011 011 101 111111 111 111 xxxxxx xxx xxx");
        $display("42 1010111001001101011101011111110xxxxxx 1010111 001 001 101011 101 011 101011 011 101 111110 111 110 xxxxxx xxx xxx");
        $display("43 1010111001001101011101011111000xxxxxx 1010111 001 001 101011 101 011 101011 011 101 111000 111 000 xxxxxx xxx xxx");
        $display("44 1010111001001101011101011010011xxxxxx 1010111 001 001 101011 101 011 101011 011 101 010011 010 011 xxxxxx xxx xxx");
        $display("45 1010111001001101011101011101011xxxxxx 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 xxxxxx xxx xxx");
        $display("46 1010111001001101011101011101011xxxx1x 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 xxxx1x x1x xxx");
        $display("47 1010111001001101011101011101011xxx01x 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 xxx01x 01x xxx");
        $display("48 1010111001001101011101011101011xxx000 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 xxx000 000 xxx");
        $display("49 1010111001001101011101011101011xxx100 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 xxx100 100 xxx");
        $display("50 1010111001001101011101011101011xxx010 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 xxx010 010 xxx");
        $display("51 1010111001001101011101011101011111111 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 111111 111 111");
        $display("52 1010111001001101011101011101011110111 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 110111 111 110");
        $display("53 1010111001001101011101011101011000111 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 000111 111 000");
        $display("54 1010111001001101011101011101011010011 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 010011 011 010");
        $display("55 1010111001001101011101011101011101011 1010111 001 001 101011 101 011 101011 011 101 101011 101 011 101011 011 101");
        #55;
    end
endmodule
module top;
endmodule
