// pattern: decl_const_var_uninit\.sv:3:16: Parse error: const declaration is missing initialization
module top;
    const var x;
endmodule
