module top;
    wire x;
    assign x = 1'bx;
endmodule
