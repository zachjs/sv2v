module top;
    initial begin
        $display("good");
        $display("good");
    end
endmodule
