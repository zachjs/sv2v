module top;
    trireg (small) x;
    trireg (medium) y;
    trireg (large) z;
endmodule
