module top;
    localparam P = 32'd1;
    localparam Q = 32'd3;
    localparam R = 832'b0;
    initial $display(P, Q, R);
endmodule
