module Example(
    input int inp,
    output int out
);
    assign out = inp * 2;
endmodule
