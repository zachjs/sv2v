interface Interface1;
    logic x;
    modport ModportA (input x);
    modport ModportB (output x);
endinterface
interface Interface2;
    logic x;
    modport ModportA (input x);
    modport ModportB (output x);
endinterface
