
module top;
    localparam P = 32'd1;
    initial $display(P);
endmodule
