// pattern: encountered continue outside of loop
module top;
    initial continue;
endmodule
