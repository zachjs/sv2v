module top;
    initial $display(1);
endmodule
