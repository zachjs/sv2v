module top;
    task foo;
        $display("foo called");
    endtask
    initial foo;
endmodule
