// pattern: localparam type "X" has no default value
module top;
    localparam type X;
endmodule
