// pattern: run_on_decl_stmt\.sv:4:20: Parse error: unexpected token in declaration
module top;
    initial begin
        integer x, byte y;
    end
endmodule
