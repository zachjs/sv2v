// pattern: unfinished conditional directive `else started at unmatched_else_end.sv:3:1
`ifdef FOO
`else
