module Module;
    Interface intf();
    assign intf.x = Package::X;
endmodule
