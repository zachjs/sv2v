module top;
    reg [5:0] a;
    wire [5:0] b;
    always @(*) a = b;
endmodule
