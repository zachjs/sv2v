module top;
    initial $display("foo");
endmodule
