module top;
endmodule
