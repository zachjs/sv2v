module top;
    Example example();
endmodule
