// pattern: unexpected keyword argument
// location: severity_task_arg.sv:4:11
module top;
    $fatal(.x("x"));
endmodule
