// pattern: missing expected `endinterface`
interface foo;
