parameter A = 1;
localparam B = A + A;
localparam C = B + B;
localparam D = C + C;
localparam E = D + D;
localparam F = E + E;
localparam G = F + F;
localparam H = G + G;
localparam I = H + H;
localparam J = I + I;
localparam K = J + J;
localparam L = K + K;
localparam M = L + L;
localparam N = M + M;
localparam O = N + N;
localparam P = O + O;
localparam Q = P + P;
localparam R = Q + Q;
localparam S = R + R;
localparam T = S + S;
localparam U = T + T;
localparam V = U + U;
localparam W = V + V;
localparam X = W + W;
localparam Y = X + X;
localparam Z = $clog2(Y + Y);
