// pattern: instantiation_not_range\.sv:3:15: Parse error: expected instantiation dimensions
module top;
    example a b();
endmodule
