// pattern: instantiation_not_ports\.sv:3:15: Parse error: expected port connections
module top;
    example a b, c();
endmodule
