// pattern: element "yes" has mismatched end label "no"
package yes;
endpackage : no
