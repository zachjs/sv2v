// pattern: declared ports w, z are not in the port list of top
module top(x, y);
    output w, x, y, z;
endmodule
