module top;
    localparam X = 5;
    localparam Y = 2;
    localparam Z = 4;
    initial $display(X, Y, Z);
endmodule
