module top;
    typedef logic T;
    T x;
    assign x = 1;
endmodule
