// pattern: encountered break outside of loop
module top;
    initial break;
endmodule
