module top;
    wire a;
    wire [1:0] b;
    wire [2:0] c;
endmodule
