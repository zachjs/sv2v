`define SIZE 4
`define NAME op
module t`NAME;
    initial $display(`SIZE'ha);
endmodule
