module top;
    wire P_T;
    assign P_T = 0;
    initial $display("%b", P_T);
endmodule
