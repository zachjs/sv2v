// pattern: bad default_nettype: "invalid"
`default_nettype invalid
module top;
    assign foo = 0;
endmodule
