// pattern: element "yes" has mismatched end label "no"
module yes;
endmodule : no
