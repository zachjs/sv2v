module top;
    logic y;
endmodule
