// pattern: missing expected `end`
module top;
    initial
        begin
            $display("FOO");
            $display("BAR");
endmodule
