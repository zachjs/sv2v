// pattern: expected typename, but found net identifier "w"
// location: typedef_not_type_net.sv:5:5
module top;
    wire w;
    w x;
endmodule
