`define ALWAYS(trigger) always @(trigger, start)
`include "always_prefix.vh"
