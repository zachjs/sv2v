package Package;
    localparam X = 1;
endpackage
