module top;
    ExampleA a();
    ExampleB b();
endmodule
