module top;
    final $display("bye");
endmodule
