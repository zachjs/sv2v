// pattern: decl_ranged_implicit\.sv:3:5: Parse error: declaration missing type information
module top;
    [1:0] x;
endmodule
