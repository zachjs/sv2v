module top;
    initial $display("%0d %0d", 1, 1);
endmodule
