module top;
    reg [5:0] s;
    initial s = 1'sb1;
endmodule
