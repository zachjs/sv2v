module top;
    wire [2:0] test;
    assign test = 3'd0;
    initial $display(test);
endmodule
