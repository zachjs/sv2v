module top;
    Example e(5'b00000);
endmodule
