// pattern: block_start_3\.sv:4:9: Parse error: expected primary token or type
module top;
    initial begin
        P::Q = 1;
    end
endmodule
