// pattern: unexpected packed range\(s\) applied to byte
module top;
    byte [1:0] x;
endmodule
