// pattern: decl_wire_var\.sv:3:10: Parse error: unexpected var after net type
module top;
    wire var x;
endmodule
