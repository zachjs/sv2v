`define ALWAYS(trigger) always_comb
`include "always_prefix.vh"
