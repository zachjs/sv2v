$display("via include: ", `__FILE__, `__LINE__);
