task fun;
endtask
function fun;
endfunction
package pop;
endpackage
module top;
endmodule
