function Function;
    input integer inp;
    return inp * 2;
endfunction
