// pattern: expected an integral number, but found 'x
module top;
    enum {
        A['x]
    } x;
endmodule
