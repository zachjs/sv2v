// pattern: size cast width 0 is not a positive integer
module top;
    initial $display((0)'(2));
endmodule
