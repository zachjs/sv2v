// pattern: instantiation_no_module\.sv:3:5: Parse error: expected module or interface name at beginning of instantiation list
module top;
    , ();
endmodule
