module top (dat_i, dat_o);
    input wire [16:0] dat_i;
    output wire [1:0] dat_o;
endmodule
