module top;
    wire x, y;
    assign y = 1;
    assign x = ~y;
endmodule
