module top;
    initial $display("hi");
endmodule
