module mod(output reg x, output wire y);
    initial x = 1;
    assign y = 1;
endmodule
