module top;
    initial $display("p %0d %b", 32, 32'bx);
    initial $display("q %0d %b", 32, 32'bx);
endmodule
