module top;
    shortreal v [2];
    real w [2];
    realtime x [2];
    string y [2];
    event z [2];
endmodule
