module top;
    initial begin
        $display(1, 2);
        $display(3, 4);
        $display(5, 5);
    end
endmodule
