// pattern: instantiation_no_label\.sv:3:13: Parse error: expected instantiation name
module top;
    example ();
endmodule
