module Example(
    input wire inp,
    output wire out
);
    assign out = ~inp;
endmodule
