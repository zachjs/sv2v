    localparam SVO_HOR_PIXELS =
        SVO_MODE == "768x576" ? 768 :
        SVO_MODE == "1280x854R" ? 1280 :
        SVO_MODE == "2560x2048R" ? 2560 :
        SVO_MODE == "1920x1200" ? 1920 :
        SVO_MODE == "480x320R" ? 480 :
        SVO_MODE == "1280x768R" ? 1280 :
        SVO_MODE == "2560x1440R" ? 2560 :
        SVO_MODE == "2048x1536" ? 2048 :
        SVO_MODE == "1024x576" ? 1024 :
        SVO_MODE == "320x200" ? 320 :
        SVO_MODE == "384x288R" ? 384 :
        SVO_MODE == "1280x1024R" ? 1280 :
        SVO_MODE == "768x576R" ? 768 :
        SVO_MODE == "2048x1536R" ? 2048 :
        SVO_MODE == "1024x576R" ? 1024 :
        SVO_MODE == "1680x1050R" ? 1680 :
        SVO_MODE == "1280x854" ? 1280 :
        SVO_MODE == "2560x2048" ? 2560 :
        SVO_MODE == "1440x900R" ? 1440 :
        SVO_MODE == "2048x1080" ? 2048 :
        SVO_MODE == "1152x768R" ? 1152 :
        SVO_MODE == "4096x2160" ? 4096 :
        SVO_MODE == "4096x2160R" ? 4096 :
        SVO_MODE == "800x480" ? 800 :
        SVO_MODE == "2560x1080R" ? 2560 :
        SVO_MODE == "1440x1080R" ? 1440 :
        SVO_MODE == "854x480" ? 854 :
        SVO_MODE == "640x480" ? 640 :
        SVO_MODE == "480x320" ? 480 :
        SVO_MODE == "1920x1200R" ? 1920 :
        SVO_MODE == "3840x2160" ? 3840 :
        SVO_MODE == "1400x1050" ? 1400 :
        SVO_MODE == "854x480R" ? 854 :
        SVO_MODE == "1680x1050" ? 1680 :
        SVO_MODE == "320x200R" ? 320 :
        SVO_MODE == "1920x1080R" ? 1920 :
        SVO_MODE == "1920x1080" ? 1920 :
        SVO_MODE == "2560x1440" ? 2560 :
        SVO_MODE == "1440x900" ? 1440 :
        SVO_MODE == "1024x600" ? 1024 :
        SVO_MODE == "1400x1050R" ? 1400 :
        SVO_MODE == "1366x768" ? 1366 :
        SVO_MODE == "1440x1080" ? 1440 :
        SVO_MODE == "1600x900" ? 1600 :
        SVO_MODE == "64x48T" ? 64 :
        SVO_MODE == "640x480R" ? 640 :
        SVO_MODE == "352x288R" ? 352 :
        SVO_MODE == "1024x768" ? 1024 :
        SVO_MODE == "800x600" ? 800 :
        SVO_MODE == "1280x960" ? 1280 :
        SVO_MODE == "1024x768R" ? 1024 :
        SVO_MODE == "1280x960R" ? 1280 :
        SVO_MODE == "1600x900R" ? 1600 :
        SVO_MODE == "800x600R" ? 800 :
        SVO_MODE == "1280x800" ? 1280 :
        SVO_MODE == "384x288" ? 384 :
        SVO_MODE == "352x288" ? 352 :
        SVO_MODE == "800x480R" ? 800 :
        SVO_MODE == "1440x960" ? 1440 :
        SVO_MODE == "3840x2160R" ? 3840 :
        SVO_MODE == "2048x1080R" ? 2048 :
        SVO_MODE == "1280x800R" ? 1280 :
        SVO_MODE == "1366x768R" ? 1366 :
        SVO_MODE == "1600x1200R" ? 1600 :
        SVO_MODE == "2560x1600" ? 2560 :
        SVO_MODE == "1600x1200" ? 1600 :
        SVO_MODE == "320x240" ? 320 :
        SVO_MODE == "1152x864" ? 1152 :
        SVO_MODE == "1440x960R" ? 1440 :
        SVO_MODE == "2560x1080" ? 2560 :
        SVO_MODE == "1152x768" ? 1152 :
        SVO_MODE == "1280x720" ? 1280 :
        SVO_MODE == "1152x864R" ? 1152 :
        SVO_MODE == "1024x600R" ? 1024 :
        SVO_MODE == "1280x1024" ? 1280 :
        SVO_MODE == "1280x768" ? 1280 :
        SVO_MODE == "1280x720R" ? 1280 :
        SVO_MODE == "2560x1600R" ? 2560 :
        SVO_MODE == "320x240R" ? 320 :
        'bx;
