// pattern: could not find package "PackageThatDoesNotExist"
module top;
    import PackageThatDoesNotExist::*;
endmodule
