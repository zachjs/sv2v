`endif
