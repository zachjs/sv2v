module top;
    initial do
        $display("hi");
    while (0);
endmodule
