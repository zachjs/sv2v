module top;
    initial $display(1);
    initial $display(8);
    initial $display(3);
endmodule
