module top;
    initial repeat (16) $display("%0d", 64);
endmodule
