// pattern: auto_dim_int\.sv:3:15: Parse error: expected comma or end of declarations
module top;
    integer x [] = 1;
endmodule
