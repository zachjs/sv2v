module top;
    reg [1:0] a[1:0];
    reg [1:0] b[1:0];

    reg [1:0] c[1:0], d[1:0];
    reg [1:0] e[1:0], f[1:0], g;
    reg [1:0] h, i[1:0];
    reg [1:0] j;

    reg [1:0] k;
endmodule
