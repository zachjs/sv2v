// pattern: decl_missing_comma\.sv:3:15: Parse error: expected comma or end of declarations
module top;
    integer a b;
endmodule
