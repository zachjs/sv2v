// pattern: Parse error: unexpected token '`'
module top;
    ``
endmodule
