module top;

    initial begin
        $display(1);
        $display(2);
        $display(3);
    end

    initial begin
        $display(1);
        $display(2);
        $display(3);
    end

    initial begin
        $display(1);
        $display(2);
        $display(3);
    end

    initial begin
        $display(1);
        $display(2);
        $display(3);
    end

endmodule
