module top;
    wire [31:0] x;
    assign x[7:0] = 1'sb1;
endmodule
