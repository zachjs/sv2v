module top;
    initial begin
        $display($signed(1'b1));
        $display($unsigned(1'sb1));
        $display($signed(1));
        $display($unsigned(1));
        $display($signed(-1));
        $display($unsigned(-1));
    end
endmodule
