module top;
    initial #1 $display("%b", 2'b11);
endmodule
