// pattern: implicit declaration of "foo" but default_nettype is none
`default_nettype none
module top;
    assign foo = 0;
endmodule
