// pattern: run_on_decl_item.sv:3:16: Parse error: unexpected comma-separated declarations
module top;
    integer x, byte y;
endmodule
