// pattern: elab_task_stray_after_args\.sv:3:12: Parse error: unexpected token after elaboration system task
module top;
    $info(), ;
endmodule
