`line 0 "asd" 3
