// pattern: instantiation_trailing_comma\.sv:3:18: Parse error: expected instantiation before ';'
module top;
    example a(), ;
endmodule
