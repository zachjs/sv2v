`define TYPE string
`include "string_type.vh"
