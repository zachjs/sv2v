// pattern: block has only end label "no"
module top;
    initial begin
        $display("Hi!");
    end : no
endmodule
