`line 1 "asd" B
