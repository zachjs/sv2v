// pattern: bad char after argument name: '#'
`define MACRO(a#)
