// pattern: element "yes" has mismatched end label "no"
interface yes;
endinterface : no
