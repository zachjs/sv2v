module top;
    wrap wrap();
endmodule
