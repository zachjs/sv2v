// pattern: block_start_2\.sv:4:9: Parse error: expected primary token or type
module top;
    initial begin
        = 1;
    end
endmodule
