module top;
    task t;
        input x;
        begin : y
            reg z;
        end
    endtask
    initial t(0);
endmodule
