module top; endmodule
`define MODULE(str) module str; initial $display(`"hello str`"); endmodule
`MODULE(example1)
`MODULE(example2)
`MODULE(example3)
`MODULE(example4)
`MODULE(example5)
`MODULE(example6)
