module top;
    /*test*/
    /*/test*/
    /*test/*/
    /*/test/*/
    initial $display("foo"/*/,"bar"/*/);
endmodule
