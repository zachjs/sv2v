// pattern: unexpected signed applied to enum
module top;
    enum {
        A, B
    } signed x;
endmodule
