// pattern: instantiation_extra_comma\.sv:3:18: Parse error: expected instantiation before ','
module top;
    example a(), , b();
endmodule
