// pattern: unfinished conditional directive `ifndef FOO started at unmatched_ifndef.sv:2:1
`ifndef FOO
