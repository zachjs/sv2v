`SOMETHING
module top;
endmodule
