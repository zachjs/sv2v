// pattern: illegal macro name: define
`define define
