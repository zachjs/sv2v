// pattern: unfinished conditional directive `ifdef FOO started at unmatched_ifdef.sv:2:1
`ifdef FOO
