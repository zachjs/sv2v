// pattern: missing expected `endinterface`
interface foo;
module bar;
endmodule
