// pattern: couldn't resolve typename "T"
// location: typedef_missing.sv:4:5
module top;
    T x;
endmodule
