// pattern: parameter_list_not_type\.sv:2:31: Parse error: unexpected non-type parameter assignment
module top #(parameter type X = 1); endmodule
