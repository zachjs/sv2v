// pattern: elab_task_stray_no_args\.sv:3:11: Parse error: unexpected token after elaboration system task
module top;
    $info , ;
endmodule
