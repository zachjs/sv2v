// pattern: Parse error
module top;
    /``* some awful garbage *``/
endmodule
