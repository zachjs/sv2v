module top;
    initial begin
        $display("Hi!");
    end//comment
endmodule
