module top;
    localparam P_X = 10;
    localparam Y = P_X;
    initial $display(Y);
endmodule
