// pattern: too few macro arguments given
`define MACRO(a, b)
`MACRO(x)
