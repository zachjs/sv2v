`define ALWAYS(trigger) always @(trigger)
`include "always_prefix.vh"
