// pattern: Could not find file "does_not_exist\.sv", included from "missing_include\.sv"
`include "does_not_exist.sv"
