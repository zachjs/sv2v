module two;
    logic x;
endmodule
