module top;
    localparam X = 1;
    localparam Y = 2;
    localparam Z = 3;
    initial $display(X, Y, Z);
endmodule
