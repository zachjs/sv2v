// pattern: element "yes" has mismatched end label "no"
module top;
    task yes;
    endtask : no
endmodule
