// pattern: expected typename, but found var identifier "v"
// location: typedef_not_type_var.sv:5:5
module top;
    var v;
    v x;
endmodule
