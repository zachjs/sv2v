// pattern: run_on_decl_item\.sv:3:16: Parse error: unexpected token in declaration
module top;
    integer x, byte y;
endmodule
