`define CASE(name, dims, a, b, c) \
module name(clock, in, out); \
    input wire clock, in; \
    output logic dims out; \
    initial out[0+a] = 0; \
    initial out[1+a] = 0; \
    initial out[2+a] = 0; \
    always @(posedge clock) begin \
 \
        out[2+a][4+b][1+c] = out[2+a][4+b][0+c]; \
        out[2+a][4+b][0+c] = out[2+a][3+b][1+c]; \
        out[2+a][3+b][1+c] = out[2+a][3+b][0+c]; \
        out[2+a][3+b][0+c] = out[2+a][2+b][1+c]; \
        out[2+a][2+b][1+c] = out[2+a][2+b][0+c]; \
        out[2+a][2+b][0+c] = out[2+a][1+b][1+c]; \
        out[2+a][1+b][1+c] = out[2+a][1+b][0+c]; \
        out[2+a][1+b][0+c] = out[2+a][0+b][1+c]; \
        out[2+a][0+b][1+c] = out[2+a][0+b][0+c]; \
        out[2+a][0+b][0+c] = out[1+a][4+b][1+c]; \
 \
        out[1+a][4+b][1+c] = out[1+a][4+b][0+c]; \
        out[1+a][4+b][0+c] = out[1+a][3+b][1+c]; \
        out[1+a][3+b][1+c] = out[1+a][3+b][0+c]; \
        out[1+a][3+b][0+c] = out[1+a][2+b][1+c]; \
        out[1+a][2+b][1+c] = out[1+a][2+b][0+c]; \
        out[1+a][2+b][0+c] = out[1+a][1+b][1+c]; \
        out[1+a][1+b][1+c] = out[1+a][1+b][0+c]; \
        out[1+a][1+b][0+c] = out[1+a][0+b][1+c]; \
        out[1+a][0+b][1+c] = out[1+a][0+b][0+c]; \
        out[1+a][0+b][0+c] = out[0+a][4+b][1+c]; \
 \
        out[0+a][4+b][1+c] = out[0+a][4+b][0+c]; \
        out[0+a][4+b][0+c] = out[0+a][3+b][1+c]; \
        out[0+a][3+b][1+c] = out[0+a][3+b][0+c]; \
        out[0+a][3+b][0+c] = out[0+a][2+b][1+c]; \
        out[0+a][2+b][1+c] = out[0+a][2+b][0+c]; \
        out[0+a][2+b][0+c] = out[0+a][1+b][1+c]; \
        out[0+a][1+b][1+c] = out[0+a][1+b][0+c]; \
        out[0+a][1+b][0+c] = out[0+a][0+b][1+c]; \
        out[0+a][0+b][1+c] = out[0+a][0+b][0+c]; \
        out[0+a][0+b][0+c] = in; \
 \
    end \
endmodule

`CASE(A1, [2:0][4:0][1:0], 0, 0, 0)
`CASE(A2, [0:2][0:4][1:0], 0, 0, 0)
`CASE(A3, [0:2][4:0][1:0], 0, 0, 0)
`CASE(A4, [2:0][0:4][1:0], 0, 0, 0)

`CASE(B1, [3:1][5:1][1:0], 1, 1, 0)
`CASE(B2, [1:3][1:5][1:0], 1, 1, 0)
`CASE(B3, [1:3][5:1][1:0], 1, 1, 0)
`CASE(B4, [3:1][1:5][1:0], 1, 1, 0)

`CASE(C1, [4:2][6:2][1:0], 2, 2, 0)
`CASE(C2, [2:4][2:6][1:0], 2, 2, 0)
`CASE(C3, [2:4][6:2][1:0], 2, 2, 0)
`CASE(C4, [4:2][2:6][1:0], 2, 2, 0)

`CASE(D1, [5:3][6:2][1:0], 3, 2, 0)
`CASE(D2, [3:5][2:6][1:0], 3, 2, 0)
`CASE(D3, [3:5][6:2][1:0], 3, 2, 0)
`CASE(D4, [5:3][2:6][1:0], 3, 2, 0)

`CASE(E1, [2:0][4:0][0:1], 0, 0, 0)
`CASE(E2, [0:2][0:4][0:1], 0, 0, 0)
`CASE(E3, [0:2][4:0][0:1], 0, 0, 0)
`CASE(E4, [2:0][0:4][0:1], 0, 0, 0)

`CASE(F1, [5:3][6:2][1:0], 3, 2, 0)
`CASE(F2, [3:5][2:6][1:0], 3, 2, 0)
`CASE(F3, [3:5][6:2][1:0], 3, 2, 0)
`CASE(F4, [5:3][2:6][1:0], 3, 2, 0)

`CASE(G1, [5:3][6:2][2:1], 3, 2, 1)
`CASE(G2, [3:5][2:6][2:1], 3, 2, 1)
`CASE(G3, [3:5][6:2][2:1], 3, 2, 1)
`CASE(G4, [5:3][2:6][2:1], 3, 2, 1)

`CASE(H1, [5:3][6:2][1:2], 3, 2, 1)
`CASE(H2, [3:5][2:6][1:2], 3, 2, 1)
`CASE(H3, [3:5][6:2][1:2], 3, 2, 1)
`CASE(H4, [5:3][2:6][1:2], 3, 2, 1)
