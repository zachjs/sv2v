module top;
    function void foo;
        $display("foo called");
    endfunction
    initial foo;
endmodule
