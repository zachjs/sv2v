// pattern: port_list_incomplete\.sv:2:17: Parse error: expected identifier
module top(input);
endmodule
