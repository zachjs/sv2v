module top(out);
    output [32 - 1:0] out;
    reg [31:0] out;
endmodule
