module top;
    wire x = 1;
    initial $display(x);
endmodule
