module apple;
    initial $display("apple");
endmodule
