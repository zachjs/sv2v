module top;
    parameter W = 8;
    reg [W - 1:0] x = 8'b1101_0100;
    wire [W - 1:0] y = 8'b0010_1011;
endmodule
