`define INPUTS inp1, inp2
`define OUTPUTS out1, out2, out3, out4, out5, out6, out7, out8, out9, outA, outB, outC
