module top;
    logic x;
endmodule
