// pattern: encountered return outside of task or function
module top;
    initial return;
endmodule
