task Task;
    $display("Hello!");
endtask
