// pattern: run_on_decl_stmt.sv:4:20: Parse error: unexpected comma-separated declarations
module top;
    initial begin
        integer x, byte y;
    end
endmodule
