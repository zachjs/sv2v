// pattern: unterminated string literal
"
