module top;
    wire o1, o2;
    mod m(o1, o2);
endmodule
