// pattern: block has only end label "no"
module top;
    if (1) begin
        wire x;
    end : no
endmodule
