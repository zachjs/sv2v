module top;
    initial begin
        $display("%b", 32'd1);
        $display("%b", 8'd2);
        $display("%b", 16'd3);
    end
endmodule
