interface orange;
    initial $display("orange");
endinterface
