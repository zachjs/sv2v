// pattern: too many macro arguments given
`define MACRO(a, b)
`MACRO(x, y, z)
