// pattern: instantiation_trailing_comma\.sv:3:16: Parse error: unexpected end of instantiation list
module top;
    example a(), ;
endmodule
