// pattern: var_var\.sv:3:9: Parse error: duplicate var modifier
module top;
    var var x = 1'b1;
endmodule
