// pattern: decl_binop_asgn\.sv:3:13: Parse error: unexpected binary assignment operator in declaration
module top;
    logic x += 1;
endmodule
