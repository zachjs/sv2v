module mod(output x, y);
    initial x = 1;
    assign y = 1;
endmodule
