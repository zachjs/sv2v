module top;
    initial $display("%b", { 8'd1, 16'd2, 32'd3, 8'd4 } );
endmodule
