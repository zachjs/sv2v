// pattern: element "yes" has mismatched end label "no"
class yes;
endclass : no
