module top;
    mod m1();
    mod #("foo") m2();
    mod #("bar") m3();
    mod #("foobar") m4();
endmodule
