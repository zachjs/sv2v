`define A
`undefineall
`ifndef A
module top;
    initial $display("hi");
endmodule
`endif
