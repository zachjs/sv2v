`default_nettype none
module top;
    assign foo = 0;
endmodule
