module top; endmodule
