module top;
    localparam Foo = 1;
    localparam Bar = 2;
    initial $display(Foo + Bar);
endmodule
