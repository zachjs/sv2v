module top;
    wire (highz0, highz1) x;
endmodule
