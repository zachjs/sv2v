// pattern: declaration type I.J appears to refer to an interface that isn't defined
module mod(I.J K);
endmodule
