// pattern: decl_signed_implicit\.sv:3:5: Parse error: declaration missing type information
module top;
    signed x;
endmodule
