module Example(
    input reg inp,
    output reg out
);
    assign out = ~inp;
endmodule
