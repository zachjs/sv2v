package P;
    typedef logic T;
endpackage
module three;
    P::T x;
endmodule
module two;
    logic x;
endmodule
