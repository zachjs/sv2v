// pattern: `elsif directive outside of an `if/`endif block
`elsif
