module top;
    initial begin
        $display(1'b0);
        $display(1'b0);
        $display(1'b1);
        $display(1'b0);
    end
endmodule
