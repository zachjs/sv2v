// pattern: unknown token '`'
// location: stray_escaped_vendor_comment.sv:4:6
module top;
    /``* some awful garbage *``/
endmodule
