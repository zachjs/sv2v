module top;
    wire P_T;
    assign P_T = 0;
    initial $display("%b", P_T);
    reg [1:0] P_U = 0;
endmodule
