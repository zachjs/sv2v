localparam UNUSED = 1;
