module top;
    localparam Foo = 1;
    initial $display(Foo);
endmodule
