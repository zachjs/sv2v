// pattern: instantiation_missing_ports\.sv:3:14: Parse error: expected port connections before delimiter
module top;
    example a, c();
endmodule
