module top;
    initial $display("%b", (12'hb03 - 12'hb07) + 12'hb10);
endmodule
