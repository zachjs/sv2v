module top;
    initial $display("Hi");
endmodule
