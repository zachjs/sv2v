module top;
    initial $display("p %0d %b", 32, 32'd1);
    initial $display("q %0d %b", 32, 32'd2);
endmodule
