// pattern: unknown token '`'
// location: double_backtick.sv:4:5
module top;
    ``
endmodule
