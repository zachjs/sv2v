// pattern: unterminated backtick string
`"
