module top;
    mod1           m1_a();
    mod1 #( 1,  2) m1_b();
    mod1 #( 0, -1) m1_c();
    mod1 #(-3, -4) m1_d();
    mod2           m2_a();
    mod2 #( 1,  2) m2_b();
    mod2 #( 0, -1) m2_c();
    mod2 #(-3, -4) m2_d();
endmodule
