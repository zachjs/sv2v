module top;
    logic [1:0] a [3];
    logic [1:0] b [3];
    always_comb a = b;
endmodule
