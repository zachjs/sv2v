`include '/dev/null'
