`define YUCK /``* some awful garbage *``/
module top;
    `YUCK
endmodule
