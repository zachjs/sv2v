// pattern: unfinished conditional directive `elsif BAR started at unmatched_elsif_end.sv:3:1
`ifdef FOO
`elsif BAR
