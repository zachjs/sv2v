`default_nettype trireg
module foo;
    not (x, y);
endmodule
`default_nettype uwire
module bar;
    not (a, b);
endmodule
