// pattern: expected beginning of macro arguments, but found 'a'
`define MACRO(a)
`MACRO asdf
