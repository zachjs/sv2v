// pattern: unexpected packed range\(s\) applied to string
module top;
    string [1:0] x;
endmodule
