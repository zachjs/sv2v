`undef RESULT

`ifndef INCLUDED
`define INCLUDED
`define RESULT 1
`else
`define RESULT 0
`endif
