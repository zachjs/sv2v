module top;
    localparam P_FOO = 10;
    initial begin
        $display(P_FOO);
    end
endmodule
