module top;
    integer x = 0;
    initial begin
        x++;
        $display(x);
    end
endmodule
