// pattern: block_start_4\.sv:4:11: Parse error: unexpected statement token
module top;
    initial begin
        a , ;
    end
endmodule
