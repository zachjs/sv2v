`define FANCY_SEEING_YOU 1337
package pkg;
    function automatic integer width_calc;
      	input integer a;
        return a+3;
    endfunction
endpackage
