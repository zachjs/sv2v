`define A