module top;
    localparam X = 10;
    initial $display(X);
endmodule
