module top;
    initial begin
        $display(`__FILE__, `__LINE__);
`line 101 "fake.v" 1
        $display(`__FILE__, `__LINE__);
    end
endmodule
