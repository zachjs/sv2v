// pattern: missing expected `endgenerate`
module top;
    generate
        initial $display("FOO");
endmodule
