// pattern: `else directive outside of an `if/`endif block
`else
