class Class;
    localparam X = 1;
endclass
