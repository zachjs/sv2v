// pattern: unexpected signed applied to string
module top;
    string signed x;
endmodule
