// pattern: missing expected `endmodule`
module foo;
module bar;
endmodule
