// pattern: missing expected `endmodule`
module foo;
