// pattern: decl_const_wire\.sv:3:5: Parse error: wire cannot be const
module top;
    const wire x = 1;
endmodule
