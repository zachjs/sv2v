module top;
    time t = 1s;
    initial $display(t);
endmodule
