interface Interface;
    logic x;
endinterface
