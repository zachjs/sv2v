`line