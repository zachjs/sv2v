// pattern: decl_trailing_comma\.sv:3:16: Parse error: unexpected token in declaration
module top;
    integer a, ;
endmodule
