module top;
    initial begin : block_name1
        integer i;
        i = 1;
        $display("%08d", i);
    end
    initial begin : block_name2
        integer i;
        i = 1;
        $display("%08d", i);
    end
endmodule
