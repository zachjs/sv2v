module top;
    initial $display("Hello!");
endmodule
