interface Interface;
    logic x;
endinterface

module Module;
    Interface i;
endmodule
