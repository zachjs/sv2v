module top;
    initial begin
        $display(signed'(4294967295));
        $display(unsigned'(4294967295));
        $display(signed'(-1));
        $display(unsigned'(-1));
    end
endmodule
