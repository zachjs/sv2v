// pattern: decl_non_blocking_asgn\.sv:3:13: Parse error: unexpected non-blocking assignment operator in declaration
module top;
    logic x <= 1;
endmodule
