module top;
    localparam AW = 16;
    wire [16:0] foo;
endmodule
