// pattern: expected a positive number, but found zero
module top;
    enum {
        A[0]
    } x;
endmodule
