`include "does_not_exist.sv"
