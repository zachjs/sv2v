module top;
    initial #(1 : 2 : 3) $display("hi");
endmodule
