// pattern: drive_strength_uninit\.sv:3:30: Parse error: net with drive strength declaration is missing initialization
module top;
    wire (supply0, supply1) x;
endmodule
