module top;
    Example e1();
    Example #(8) e2();
    Example #(9) e3();
endmodule
