// pattern: charge_strength_non_trireg\.sv:3:5: Parse error: only trireg can have a charge strength
module top;
    wire (small) x;
endmodule
