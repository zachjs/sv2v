// pattern: macro definition missing argument name
`define MACRO()
