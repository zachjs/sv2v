`default_nettype none
`resetall
module top;
    assign y = 1;
    assign x = ~y;
endmodule
