// pattern: invalid macro definition argument: "#"
`define MACRO(#)
