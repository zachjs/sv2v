module top;
    initial $display("Module1 P=%0d", 5);
endmodule
