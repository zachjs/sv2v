module top;
    mod #("FOO") m1();
    mod #("BAR") m2();
endmodule
