extern module foo(input x, output y);
