// pattern: Undefined macro: SOMETHING
`SOMETHING
module top;
endmodule
