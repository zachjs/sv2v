module top;
    wire [31:0] x = 1'sb1;
endmodule
