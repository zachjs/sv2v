// pattern: block_start_1\.sv:4:9: Parse error: expected primary token or type
module top;
    initial begin
        ,;
    end
endmodule
