module top;
    localparam Bar = 2;
    initial $display(Bar);
endmodule
