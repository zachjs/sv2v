module top;
    initial begin
        $display("A %0d", 32);
        $display("B %0d", 10);
        $display("C %0d", 32);
        $display("D %0d", 6);
        $display("E %0d", 32);
    end
endmodule
